----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/31/2025 06:27:35 PM
-- Design Name: 
-- Module Name: big_alu - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity big_alu is
    Generic ( WIDTH : positive := 23);
    Port ( op1 : in STD_LOGIC_VECTOR(WIDTH-1 downto 0);
           op2 : in STD_LOGIC_VECTOR(WIDTH-1 downto 0);
           sel : in STD_LOGIC;
           en : in STD_LOGIC;
           shift_flag : in STD_LOGIC;
           
           carry : out STD_LOGIC_VECTOR(1 downto 0); --carry signal koji sadrzi implicitnu vrednost - hidden value
           result : out STD_LOGIC_VECTOR(WIDTH-1 downto 0));
end big_alu;

architecture Behavioral of big_alu is

    --signal result_s ima 2 dodatna bita u odnosu na result zato sto je neophodno izracunati skrivenu vrednost
    signal result_s: unsigned(WIDTH+1 downto 0):= (others=>'0');  --uvodjenje ovog unutrasnjeg signala ce verovatno ubaciti latch kako bi memorisao stanje medjusignala?

begin

    alu: process (en, sel, op1, op2) is
    -- da li je enable signal neophodan u sensitivy listi? NARAVNO 
    begin
      if(en = '1') then
        if(sel ='0') then
            
            --result <= std_logic_vector(unsigned(op1) + unsigned(op2));
            
            --result_s <= ('0' & unsigned(op1)) + ('0' & unsigned(op2));
            
            if(shift_flag = '0') then
              result_s <= ("01"&unsigned(op1))  +  ("01"&unsigned(op2));
            else
              result_s <= ("00"&unsigned(op1))  +  ("01"&unsigned(op2));
            end if;
            
          else
            --ALWAYS SUBTRACTING OP1 FROM OP2 because OP1 is always set to smaller shifted or not shifted, always smaller
            if(shift_flag = '0') then
              --result <= std_logic_vector(unsigned(op1) + (not(unsigned(op2))+1));
              --result_s <= ('0' & unsigned(op1)) + (not('0' & unsigned(op2)) + 1);
              result_s <= ("01"&unsigned(op2))  -  ("01"&unsigned(op1));
            else
              result_s <= ("01"&unsigned(op2))  -  ("00"&unsigned(op1));
            end if;
  
        end if;
        --carry <= std_logic(result_s(WIDTH)); --uzme msb kao carry out signal
      else
        result_s <= (others => '0');
        --carry <= '0';
      end if;
      
    end process alu;
    
    --carry <= std_logic(result_s(WIDTH));
    carry <= std_logic_vector(result_s(WIDTH+1 downto WIDTH));
    result <= std_logic_vector(result_s(WIDTH-1 downto 0));

end Behavioral;
